`include "apb_interface.sv"
`include "rtl\apb_mem.sv"