import uvm_pkg::*;

class base_test extends uvm_test
    `uvm_component_utils(base_test)
    

endclass