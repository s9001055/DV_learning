`include "apb_interface.sv"